
`define Store 4'b0000    
`define INPM 4'b0001  
`define INSW 4'b0010
`define ADD 4'b0011
`define ADDI 4'b0100
`define MUL 4'b0101
`define MULI 4'b0110
`define SW80 4'b0111
`define SW81 4'b1000