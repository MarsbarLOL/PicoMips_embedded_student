//
`define RA 2'b00
`define RB 2'b01
`define RADD 2'b10
`define R_mul 2'b11


